interface dff_intf();

    logic clk;
    logic rst;
    logic din;
    logic dout;

endinterface: dff_intf
