interface mul_intf();

    logic [3:0] a;
    logic [3:0] b;
    logic [7:0] y;

endinterface: mul_intf
