class rand_baud extends uvm_sequence #(uart_transaction); 
// random baud rate 
// 1 stop bit
// parity en
// parity type : random
    `uvm_object_utils(rand_baud)

    uart_transaction trans;

    function new(string name = "rand_baud");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = rand_baud_1_stop;
            trans.length = 8;
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b1;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud

class rand_baud_two_stop extends uvm_sequence #(uart_transaction); 
// random baud rate 
// 2 stop bits
// parity en
// parity type : random
    `uvm_object_utils(rand_baud_two_stop)

    uart_transaction trans;

    function new(string name = "rand_baud_two_stop");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = rand_baud_2_stop;
            trans.length = 8;
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b1;
            trans.stop2 = 1'b1;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_two_stop

class rand_baud_len5_p extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len5_p)

    uart_transaction trans;

    function new(string name = "rand_baud_len5_p");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length5wp;
            trans.length = 5;
            trans.tx_data = {3'b000, trans.tx_data[7:3]}; // 000 5LSB - generated by PRNG
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b1;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len5_p

class rand_baud_len6_p extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len6_p)

    uart_transaction trans;

    function new(string name = "rand_baud_len6_p");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length6wp;
            trans.length = 6;
            trans.tx_data = {2'b00, trans.tx_data[7:2]}; // 000 5LSB - generated by PRNG
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b1;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len6_p

class rand_baud_len7_p extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len7_p)

    uart_transaction trans;

    function new(string name = "rand_baud_len7_p");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length7wp;
            trans.length = 7;
            trans.tx_data = {1'b0, trans.tx_data[7:2]}; // 000 5LSB - generated by PRNG
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b1;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len7_p

class rand_baud_len8_p extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len8_p)

    uart_transaction trans;

    function new(string name = "rand_baud_len8_p");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length8wp;
            trans.length = 8;
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b1;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len8_p

class rand_baud_len5_wop extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len5_wop)

    uart_transaction trans;

    function new(string name = "rand_baud_len5_wop");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length5wop;
            trans.length = 5;
            trans.tx_data = {3'b000, trans.tx_data[7:3]}; // 000 5LSB - generated by PRNG
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b0;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len5_wop

class rand_baud_len6_wop extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len6_wop)

    uart_transaction trans;

    function new(string name = "rand_baud_len6_wop");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length6wop;
            trans.length = 6;
            trans.tx_data = {2'b00, trans.tx_data[7:2]}; // 00 6LSB - generated by PRNG
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b0;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len6_wop

class rand_baud_len7_wop extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len7_wop)

    uart_transaction trans;

    function new(string name = "rand_baud_len7_wop");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length7wop;
            trans.length = 7;
            trans.tx_data = {1'b0, trans.tx_data[7:2]}; // 0 7LSB - generated by PRNG
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b0;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len7_wop

class rand_baud_len8_wop extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_baud_len8_wop)

    uart_transaction trans;

    function new(string name = "rand_baud_len8_wop");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = length8wop;
            trans.length = 8;
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b0;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_baud_len8_wop

class rand_length extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_length)

    uart_transaction trans;

    function new(string name = "rand_length");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = rand_length_1_stop;
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b0;
            trans.stop2 = 1'b0;
            finish_item(trans);
        end
    endtask:body
endclass: rand_length

class rand_length_two_stop extends uvm_sequence #(uart_transaction);
    `uvm_object_utils(rand_length_two_stop)

    uart_transaction trans;

    function new(string name = "rand_length_two_stop");
        super.new(name);
    endfunction: new

    task body();
        repeat(5) begin
            trans = uart_transaction::type_id::create("trans");
            start_item(trans); //send request to sequencer that we have new data
            assert(trans.randomize());
            trans.oper = rand_length_2_stop;
            trans.rst = 1'b0;
            trans.tx_start = 1'b1;
            trans.rx_start = 1'b1;
            trans.parity_en = 1'b0;
            trans.stop2 = 1'b1;
            finish_item(trans);
        end
    endtask:body
endclass: rand_length_two_stop
